[PathToGnuPG]
PathToGnuPG=c:/Program Files/gnu/gnupg/gpg.exe

[PresetUserInformation]
Name=�e�X�g����
ID=012345678

[PresetRecipientInformation]
Count=2
PublicKeyTitle1=�e�X�g���t��P
PublicKeyFile1=P_Test01.asc
IsRecipient1=1
PublicKeyTitle2=�e�X�g�����̂�
PublicKeyFile2=P_Test02.asc
IsRecipient2=0
